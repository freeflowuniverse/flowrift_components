module components

pub struct Accordion {

}