module contact

pub struct ContactForm {
pub:
	title       string  = 'Get in touch'
	description string  = 'This is a section of some simple filler text, also known as placeholder text. It shares some characteristics of a real written text but is random or otherwise generated.'
	post_url    string  = '/' // where the form content will be posted to
	name_inputs []Input = [
		Input{
			label: 'First name'
			id: 'first-name'
		},
		Input{
			label: 'Last name'
			id: 'last-name'
		},
	]
	contact_inputs []Input = [
		Input{
			label: 'Company'
			id: 'company'
		},
		Input{
			label: 'Email'
			id: 'email'
		},
		Input{
			label: 'Subject'
			id: 'subject'
		},
	]
	message Input = Input{
		label: 'Message'
		id: 'message'
	}
}

pub struct Input {
pub:
	label string
	id    string
}

pub fn (component ContactForm) html() string {
	return $tmpl('./templates/form.html')
}
