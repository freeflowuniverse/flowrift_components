module logos

pub struct Logos {
pub mut:
	title       string    = 'logos'
    logos    []Logo = []Logo{len: 4}
}

pub struct Logo {
pub mut:
	title       string = 'A logo'
	img   string = 'data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAAUYAAACbCAMAAAAp3sKHAAAAjVBMVEX///8AAADy8vKysrKlpaX8/Pzp6enu7u739/eurq61tbXa2tr4+Pjl5eXU1NTd3d19fX3Dw8PKyspXV1eNjY2goKBpaWkwMDBcXFy9vb1vb2+oqKiHh4dOTk4XFxeBgYE8PDxqampFRUWXl5cfHx8NDQ0tLS1BQUGMjIwWFhYdHR04ODgLCwt1dXUmJiZ2m8KFAAAOlUlEQVR4nO1dZ2OyMBB24OQVXFhnq9Jt7f//ea/ZdyEBHCjWPJ9aZnhyuZVLrFQcHBwcHBwcHBwcHBwcHBwcHBwc8qAZdKP+6IljNR8vBmH71o26J4Td5eitasa27w1bt25g+dHuTC0EQozGA8elHbVJDg453vb15q3bW06E+Unk6A8at2506VA7mkWC1cKNb4TdSTQesPZqt257eeBBYib9cRxFURx/7ier9xwy2b1180uCf4LB2ODRNA5eZDxJp7Mf3qDVpUOfcrFIH54Hl3KdMrhnV2prifFNmdgPM9VcI4hXViajR7fcippl9sWNwYuNyPHJEWN7eIg+39+qb7uJd7cuae1bMjHIdYM//jITuTyFyODzFz1kcrdivfigH/Ac577DX1ok8kgO/sU/iWd83S2PlUqr2Tyy9YORkcjFMc8YGx+xP64h946WkYXnfJrhgIFZoqvVp0nUK7LhpUPX5FGu8nEwt7FIMX2sFOfQ5APlMPntp1QWD3iwODM0JSqzRnYLyN2yb6RxfYW2lwo9Q7YyfVDKnFJ8UAAzizgG12p/aWAisp5yPXdVI/I3FuZdfynUxOeVGl8mhEn/Z2QVSMbcG4lYWt/gjl8W2Qfsv8nVGl8mBMm0pUVDdtlZwjLMuytX6ZPphSs1vGxIKjmzJ83O+RUpdxQghmI8v1yn1SVErPP4a5hoiOiZeQWx+BYmruhcq9W3gZfyfbWE95Mc2F9CGH111QpdsaXH7jbZkwv1dK2VCPH0hAdXhwfzbhv8TEg/Lt7yUuHbQA3CXuNRI71OD27hfKSmBV8tYvyXwGQoNWweajzuUPIo5tx+21hkPuj60g0vFzyThOnQvPFnGB+zvNBK+ZlzfC9Pr//xHA///Az9X9cEEly+0E5h6yISP97lW14qVPN9Zu/ZxmOAT7yi2wKmF6ubAlpeJoiwIzvE0FwfxSM+Dh3LQNyzSj7ub6HDP/Qt+9JPC18RPKrSOEEs57ZGhTS9TJDzqzmu7SIa36S9hlmM3eQljuLlBgbk87SH/g1sk4PUDuz5PMnj39U0/HXrQiA/NlfhDi6clPrUMj1L8foIFUEq9MiXm+4hikTw82pnMf9c+T1DZROG+W5oIpLYTfay1MmDVJ4ONEaygeWRJcQtJO7/dk4HoCO/OS+NMB0mHMIN+6cLTfaqc8dFJ8ciPp5GnDqjZpiN9IMarHVfRtuP1T4aPhCHFVFTSnBEZSjyt6n2IyH3+2Vb1sgu0CwPJqfQiBI+bFgH888Ly9/qnqy8KjU5qnQe+tsFFTiTR99NQkPFbP1BEOYeRsgNL6RhrJrlLiYTewM9V1it/q7mn4tB+C/jVjhlWMjYa7Bnp5VqlABhp5+yEoFgtOymJaxh4KK0YqO/sVn8f/4sWm6m2+12NZkvo/qwl95VPL9Z3qR5GJkLaw2YdmweNMxSKHEkiQ5DJsL3Nsby8tHY7mbxibTnMz+2IATWlQcW7Dyz1MA6SPlw+p+PL5yl14/uLQpZZOXG1k9p1HrBoLuIoqjrJ896P4VVsPXSUjEpX2qKjOHcgagXYF20hm/M0WuCR1xpJQN17eXNYTd+Sa7b08SazHkUpFdnHyeRSGAqtwW6VWQeebpbyka+Zd08v7HVjJV4Pkj6Dj631qegWn/ax4WsfuxYG5AHP8msIcyFM0PAratkQ59OtKCm7oW1e7Kgn4tjqJcdaAAlNCzsL2BQD5/T25CNZNEDOMmIE97kSOMhHaxQZQIfxJosLuDlpfaFeRxyEPBkHmqs3/VmZ2ftMjoyFxKdC6YK1/SAyFn8oP8y8It6ANinhryE/Z/0cTX88Bv5El6gDGq8R6fnhenmdeqvuxHQltPVLiWJTaAX20I1QV1HuZCbnrasoJNvf3/arqZLHkpuxGEwQymV70Cj1YYO+lrV7WBYnOOGIhZ/J+PO0G8xl1npN24lDj5EN96bFbledAwjQtpm6QeQTg/0299H82XcmQ2DsJkQira6TMXRckKX16fppUQJsLkhPvLW4jE+2kPn9ASK/LrdS93Hj1ECpU3I14bePiGcmisOxYPaSWmXe/Ct1bf+IitkgYItUx1KK/ADiZ7RQPtZlAgLYYzwNSevvOMOWN+USVX7KZjmktvaKuFIOw9OUY9ICjEx62IIPOfJByPzIWRVTfFIhdlNszP9NrhJDJ2NftWpdsYzMQDPsTZY7g5ADKKParDil/aC9AbIZ4u/8yzjwGpPDgz5PNh6dd3P69NqNOkvY68+G/qcfBHnckWepP3URArRFTYXSiVq7DFXTwYMeg0J0Lkj9IU+ZOYpGvYyLKRm1IUHKHsQ9J8co2apEk/irrdBeE8t+p2TUlgLlA1L6yTD11AAGokEKTvhJ+3q77Qfdwa+OdOhx6hclNRYSbbFUhaEz2IWp+/as47CQeK+bOdU+y2jnkJIhU41yIETI6mmsMmgTq5P51jP45nmd+g5O16OoUyzNFCSWXPALGSVST8KRX97XG+eOOtLJpZtiX41o5Wy/FwKlu50gUYSA6hmXomJyciCTLoN44MY9DICP3GleUzzk0wroBZM5YcYskG5MLK+FfSXPR0y+wItgYDFEkS1KuEhNDYy0sIHqyY0pp849YNYUZGoZMas4bgw7ug/KIlA9VH7LBrpYDMreRXPWWhsAZdHfwR0h0n/q0VdTGxnmVEwtyUyCFA3MP0hPSg6VvzYtML4aaNyEvwQNaiob6aKiJNpZArFqBJUMGjOKkETmrD2MPVA2qa6X8h+YxjtV1YlWRVTVlLGutojpKkmrJpXaRPUcGupw9SGFzDxNGeVjwAVOlOBnPL8MmlMvh3OspL/VbygqZB/PX/Y9cb7Ed5ahoBKkpzTCJXxp/IjO4rQbWVRNo2PLapYUQDMLZRXtfGQE0/y8RjqTZYcZ4+PK4MTDUMzKgDKCYXDvzeLxuPYmwX0YC2o4129GrAV8KHDCrDL/UoajXycCFNI/kaii2k+I8vDRDw52ZRJ44GGeuwZ4zk4L0bdJWUZZS6ojXKOH8sZS9EOVeKuo/amo4sYpLb+rgClSWi0mywuX1w3Lyva2lv52YrlU8G0q+4//1PvOjrjjvIEVPEqCRA0wi0QOZ4iNuKF6E6BMSBOs0obRUCnEBq1HAMAd534+wdaEaZ0MFgy/rxFEaytz1gxgI02jqYR5n8+4GcoGi1TglNKuugGIDo0+6Kch5qikehGXFgJIOJYHrS2sNZWoQcL0c8sTuDuCXoKcAqOpRHl09nNG0AAgV18qJLgrLeVTl3iNr0oGglTqs9H0aJ+wMKr12eBMmf8rLaCR8YMPHt+7gwN5/E1SBw6gUZMETumfHkwSeX1wk5yix5ynqvNpuoR1sXKeazJ9nmoseZwjo/kX9w2qRhFLxz3nQaIYTSVHQg08XGTuljpcf9XCQF9AbUPLPwYaBlgUgoh7GqobFWEmnkYjxvxFwlmZS9ZtBsX4y1S2upa7mxdoOBIapeXWoKNo2jE67W++VFFIxUXMlZlzFaHRD4dzrd+5bXSm+TdYZjCCOCYtgwcLq3YN5XezVY/cAZqMnXIiATuyBE0/tOCPKEllAdE9REZWzt1V9hZblbb7bTvHcxcQ/mYbeV1cX4McwU16E5ZplNMUzXiq2SAf6FKPyUx8xDZifw04iVvYHZD0RjKzzLmvn3oHAPnVeShkrt7VcBVtkWiyQSHzLOqjskqOMwLoH+3Q+BB56Ux0L3gb3lKo5F9+Le2LWttsEQzdSsQ/QovH6+9qVJ/Vx2TKb3msB6/bCYrPv/R0u8Stqi9T957Ngydlp9Gw356iiWdRjk/v9rH0cFBieK9aWrEkFXU66cWMLrvVdrhIJoD8/9qWZ1DHcomeJh1FuAUGOuTctBY8wz1AMB9UmOR+2qZGUd6qaJR9og+A9GC1tDQiK32foZnUsqJyr8uu7bBVBaSVQjfXBizhzDa1hweLVllxge8SikurH8JS4mNlRDoC/XqlA+9xfmX/uRDIxmm/cw71kRcWN9bkoYoJFAqSPBRyyhAYQ+Q/4BnIQaI85leV0XFP6vXCliQHCRTfwe8b+L60G/ykLjW9A9KfGPfJvQLWw/lkshDjYwEODXkgms4MQCSJsxrskeW6oXpBV/FrGowZF+OhJ4vkk9cg4OpZZUspBC6GlUcgAIh2lm6m4XAR2tqcUpRWww0jq0C15AoeJRfgfhoWKcI+1yFCp2GrZz0KJjisOZ3qmn+pkKBGzW0jCM7H0xVFuKcRnDDM+iFqZpgFXZZs6M1qsDlimxrneuXSP6l/WZTjk2OT8fJ1aMvRtehyWNNw5nOXPkpu7mHs1VswBqqiJpgZtymHFV/pghjsT+Ck7OsWEds3Z017MSRdUu3ph8EQc90r7+c7DOXHhqbArYPsA/7XcHL408pq5/cauc7gwGZwDoO6/KbwrffBEmRfIs9NrMbLjfX94h9QUJm2fBifYVVhyCan1XSfoSHYBqdPlF+GfjAm5/qSgApqHm0J0m5Zfc6W4aoFzOlH87Ghh/a2u6jkvw45my//vn62ESGCRXU4iu3ViX+4FFS5TCYdbvdwSAIy8FfJpB7fu090aR1sxfb3glQNunSOYhM8MTJ3W/fi7ydn+zrLw1SPfd1P3tj2IAm2dIqhx3SgAzMHe08Uy4g1/xRf3vhfKBk1d/eYLxIoDF968bcLdBs513s3VNKoPmux/utqUth7cb0BQDnvx7yF7suAzTvfus01P3i043pSwAWRNrWhTtkAgrj1ZM7fwY9N6YvAWhh/v6PWBQGWEn2CL+/UBDgZNYj/ABDQYBFQrduyx0D0OhSjacDeN9u+uB0gEpNl905HUOnGi8BleBhe0FWZt2H+YWVS0IWNtIy6sY4GNQdj8dDzgvS2o9Fa1Gr/PHfwi4GYn0YLapd9FqVSsl/BKCcEAWGNIapdbxO6BI9p6ADDXXQ6RZb6/130ZcWxuEcfDrn+yLo2ZdAODg4ODg4ODg4ODg4ODg4OJQa/wGfU6xbqlrh8QAAAABJRU5ErkJggg=='

}

pub fn (component Logos) html() string {
	return $tmpl('./templates/logos.html')
}
