module reviews

import freeflowuniverse.crystallib.data.ourtime

pub struct NewsLetter {
pub:
	description        string
	signup       string
	legal string
	terms_conditions_link string
	image   string [required]
}
