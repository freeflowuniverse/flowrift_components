module cta

import freeflowuniverse.crystallib.core.playbook
// import freeflowuniverse.crystallib.data.ourtime
// import freeflowuniverse.webcomponents.components.stars

const actor = 'flowrift'

pub fn process(txt string) !string {
	mut plbook := playbook.new(text: txt)!

	if plbook.action_exists_once(actor: cta.actor, name: 'cta') {
		a := plbook.action_get_by_name(actor: cta.actor, name: 'cta')!
		mut d := a.params.decode[CTA]()!
		return process_from_model(d)!
	}

	return ''
}

pub fn process_from_model(component CTA) !string {
	return component.html()
}
