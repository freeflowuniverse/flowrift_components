module components

import veb

// @['/slides/:name']
// pub fn (app &App) slides(mut ctx Context, name string) veb.Result {
// 	doc := model_web_example()
// 	// d := $tmpl('templates/index.html')
// 	panic('implement')
// 	// return ctx.html(d)
// }
